module DATA_SYNC #(
    parameter NUM_STAGES = 2,        // Number of flip-flop stages for synchronization
    parameter BUS_WIDTH = 8          // Width of the bus (number of bits in Unsync_bus and sync_bus)
) (
    input  wire                 CLK,         // Destination domain clock
    input  wire                 RST,         // Active-low asynchronous reset
    input  wire [BUS_WIDTH-1:0] unsync_bus,  // Unsynchronized input bus
    input  wire                 bus_enable,  // Enable signal from the source clock domain
    output reg  [BUS_WIDTH-1:0] sync_bus,    // Synchronized output bus after synchronization
    output reg                  enable_pulse // Synchronized enable pulse, generated based on bus_enable
);

reg [NUM_STAGES - 1 : 0] sync_reg;  // Multi-stage flip-flop register chain to synchronize the bus_enable signal
reg in_flop;                        // A flip-flop used for pulse generation

wire pulse_ou;                      // Output pulse signal generated by detecting transitions in bus_enable
wire unsync_reg;                    // Intermediate signal for unsynchronized data (not used in this code, can be removed)

// Multi-stage synchronization
always @(posedge CLK, negedge RST) 
begin
    if(!RST)
        begin
            sync_reg <= 'b0;
        end
    else
        begin
            sync_reg <= {sync_reg[NUM_STAGES - 2 : 0], bus_enable}; // Shift the bus_enable signal through the flip-flops
        end
end

// Capture the final flip-flop stage output
always @(posedge CLK, negedge RST) 
begin
    if(!RST)
        begin
            in_flop <= 1'b0;
        end
    else
        begin
            in_flop <= sync_reg[NUM_STAGES - 1]; // Capture the last flip-flop output from sync_reg
        end
end

// Pulse generation: Detect a rising edge by comparing the last two stages of sync_reg
assign pulse_ou = sync_reg[NUM_STAGES - 1] & (~in_flop);

// Update the synchronized bus
always @(posedge CLK, negedge RST) 
begin
    if(!RST)
        begin
            sync_bus <= 'b0;
        end
    else if (pulse_ou)
        begin
            sync_bus <= unsync_bus;  // Update the synchronized bus with the unsynchronized bus data when pulse_ou is high
        end
end

// Update the enable_pulse signal with the generated pulse_ou
always @(posedge CLK, negedge RST) 
begin
    if(!RST)
        begin
            enable_pulse <= 1'b0;
        end
    else
        begin
            enable_pulse <= pulse_ou; // Set enable_pulse when pulse_ou is high
        end
end

endmodule
